module SimpleModule (
    input  logic port1,
    output logic port2
);

    assign port1 = port2;

endmodule : SimpleModule
